`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.06.2023 21:16:12
// Design Name: 
// Module Name: user_interface
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module user_interface(
    input clk,
    output [3:0] delay,
    output [3:0] mode,
    output [3:0] threshold,
    output [3:0] corner_freq,
    output [3:0] amplitude_scale,
    output [3:0] time_scale
    );
endmodule
