`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.07.2023 09:31:41
// Design Name: 
// Module Name: trigger_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module trigger_rom(
    input logic clk,
    input logic data,
    output logic data_output_trigger,
    output logic data_output_display,
    output logic delay
    );
endmodule
